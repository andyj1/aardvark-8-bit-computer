//////////////////////////////////////////////////////////////////////////////////
//
// School: The Cooper Union
// Course: ECE151A Spring 2016
// Assignment: Final Project -- 8-bit computer
// Group members: Andy Jeong, Brenda So, Gordon Macshane
// Date: 04/20/2016
// DUT (Device Under Testing)
//////////////////////////////////////////////////////////////////////////////////
module main_tb();

//?????????????Input Ports?????????????????????????????
// inputs to the DUT are reg type
reg [4:0]data1;

//?????????????Output Ports????????????????????????????
// outputs from the DUT are wire type
wire [7:0]result;

//??????----?-??????Instructions---???????????????--???

// instantiate the DUT using named instantiation
signext5 signext(result, data1);

//initial blocks are sequential and start at time 0
initial
begin
	$display("<<Starting the Simulation>>");
	data1 = 5'b10101;
	$display("data1: %b result: %b", data1, result);
	$display("data1: %d result: %d", data1, result);
end

endmodule
		