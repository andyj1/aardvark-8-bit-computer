//////////////////////////////////////////////////////////////////////////////////
// Created by: Team Aardvark
// Course: Cooper Union ECE151A Spring 2016
// Professor: Professor Marano
// Module Name: 
// Description: 
//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ns

module register_file ();

//-------------Input-------------------
input t0;	//slt_0 register 
input t1;	//slt_1 register 
//-------------Output------------------
output [2:0] ALUctrlbits;

//-------------Input ports Data Type-------------------
wire t0;	
wire t1;

//-------------Output Ports Data Type------------------


//------------------Instructions-----------------------


endmodule
